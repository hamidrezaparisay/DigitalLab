module ins_memory(ins_address,ins,clk);
input clk;
input [9:0] ins_address;
output [31:0] ins;
reg [31:0] ins_reg;
reg [7:0] a [1024:0];

assign ins[31:24]=a[ins_address];
assign ins[23:16]=a[ins_address+1];
assign ins[15:8]=a[ins_address+2];
assign ins[7:0]=a[ins_address+3];

initial begin
	a[0]=8'b00000001;
	a[1]=8'b01000000;
	a[2]=8'b00000101;
	a[3]=8'b00010011;

	a[4]=8'b00000000;
	a[5]=8'b00010000;
	a[6]=8'b00000101;
	a[7]=8'b10010011;

	a[8]=8'b00000000;
	a[9]=8'b00000000;
	a[10]=8'b00000110;
	a[11]=8'b00010011;

	a[12]=8'b00000000;
	a[13]=8'b10100101;
	a[14]=8'b10000100;
	a[15]=8'b01100011;

	a[16]=8'b00000000;
	a[17]=8'b10110110;
	a[18]=8'b00000110;
	a[19]=8'b00110011;

	a[20]=8'b00000000;
	a[21]=8'b00010101;
	a[22]=8'b10000101;
	a[23]=8'b10010011;

	a[24]=8'b11111110;
	a[25]=8'b00000000;
	a[26]=8'b00001101;
	a[27]=8'b11100011;

	a[28]=8'b00000000;
	a[29]=8'b11000000;
	a[30]=8'b00110000;
	a[31]=8'b00100011;
		
end
endmodule